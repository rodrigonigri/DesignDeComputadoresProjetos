library ieee;
use ieee.std_logic_1164.all;

entity UnidadeControleULA is
  port ( opcode : in std_logic_vector(5 downto 0);
			tipoR : in std_logic;
			funct : in std_logic_vector(5 downto 0);
         operacao : out std_logic
  );
end entity;

architecture comportamento of UnidadeControleULA is

  constant lw  : std_logic_vector(5 downto 0) := "100011";
  constant sw  : std_logic_vector(5 downto 0) := "101011";
  constant beq : std_logic_vector(5 downto 0) := "000100";
  constant jmp : std_logic_vector(5 downto 0) := "000010";
  constant op_r : std_logic_vector(5 downto 0) := "000000"; 
  constant funct_add : std_logic_vector(5 downto 0) := "100000";
  constant funct_sub : std_logic_vector(5 downto 0) := "100010";
  

  begin
  -- seletor da operação = "1" quando soma e "0" quando subtração
  -- soma quando:
  	-- tipoR = "0" e opcode = lw
	-- tipoR = "0" e opcode = sw
	-- tipoR = "1" e funct = add
  -- subtracao quando:
	-- tipoR = "0" e opcode = beq
	-- tipoR = "1" e funct = sub

  
  operacao <= '1' when tipoR = '0' and opcode = lw else 
				  '1' when tipoR = '0' and opcode = sw else 
				  '1' when tipoR = '1' and funct = funct_add else 
				  '0' when tipoR = '0' and opcode = beq else 
				  '0' when tipoR = '1' and funct = funct_sub else 
				  '0';
  
			  
end architecture;